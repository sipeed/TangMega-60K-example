`define MODULE_NAME SerDes_Top
