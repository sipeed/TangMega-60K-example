`define module_name PCIE_Controller_Top
`define tl_clk_freq 100
`define msi_int
