parameter DRP_NUM = 4;
